
`ifndef _MATRIX_H_
`define _MATRIX_H_

  `define MAX_VALUE 16
  `define NUM_X     4
  `define NUM_Y     4

`endif
